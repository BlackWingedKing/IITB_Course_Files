Q4(3)
*Passive Components
R 1 2 1k
C 2 0 100n

*ac source of 10Vpp
vin 1 0 dc 0 ac 5

*vary frequency from 50-50khz
.ac dec 10 50 50k

.control
run

*plot the outputs
plot vdb(2) xlog
plot {57.29*vp(2)} xlog
*v(2) is output voltage and v(1) is input voltage

.endc
.end
