library ieee;
use ieee.std_logic_1164.all;

entity  dflip is
  port(D, CLK, RST : in std_logic; 
		Q, Qbar : out std_logic);
end entity;
architecture behave of dflip is
begin 
   process (CLK,RST) 
   begin
		if (RST = '1') then
			Q <= '0';
			Qbar <= '1';
		elsif CLK'event and (CLK = '1') then
			Q <= D;
			Qbar <= not D;
		end if;
   end process;
end behave;