Q4(3) Scmidtt Trigger
.include ua741.txt
x1 1 2 3 4 5 UA741
R1 0 1 6.8k
R2 1 5 10K
Vin 2 0 sin(0 10 1kHz)
Vss 3 0 dc 12
Vdd 0 4 dc 12

.tran 0.001ms 5ms

.control
run

plot v(5) vs v(2)
plot v(5) v(2)
.endc
.end
