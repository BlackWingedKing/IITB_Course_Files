Lab5 light condition Q1
.include Solar_Cell8.txt

*define the Cell and others 
xs 1 0 solar_cell
vi 1 0 dc 0 ac 0


*analysis
.dc temp 35 75 5

.control
run

*plot the required graphs
plot i(vi)
.endc
.end
