Q6
.include bc547.txt
*after solving Rc=3k,Re=2k,R1=27k given R2=10k
*passive elements in the cicuit
Re 0 1 2k
R2 0 2 10k
Rc 6 7 3k
R1 2 7 27k

Rl 9 0 1k

Cc 5 9 50u
Ce 1 0 50u
Cb 2 8 50u

*biasing voltage
Vba 7 0 dc 10v

*voltage sources for measuring currents
vie 3 1 dc 0v
vic 6 5 dc 0v
vib 2 4 dc 0v

*nodes of the transistor
q1 5 4 3 bc547a
*input voltage 
vin 8 0 dc 0 ac 10

*transient analysis
.ac dec 10 10Hz 100KHz

.control
run
plot v(9)
.endc
.end
