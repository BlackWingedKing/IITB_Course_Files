Lab3 Question1
.include Diode_1N914.txt
.include red_5mm.txt
.include green_5mm.txt
.include blue_5mm.txt
.include yellow_5mm.txt
.include white_5mm.txt

*defining the diode
d1 1 2 1N914
dr 1 3 RED
db 1 4 BLUE
dy 1 5 YELLOW
dg 1 6 GREEN
dw 1 7 WHITE

*Current sources for measuring current across diode
v1 2 8 dc 0 ac 0
vr 3 9 dc 0 ac 0
vb 4 10 dc 0 ac 0
vy 5 11 dc 0 ac 0
vg 6 12 dc 0 ac 0
vw 7 13 dc 0 ac 0

*Resistance measurement
r1 8 0 100
rr 9 0 100
rb 10 0 100
ry 11 0 100
rg 12 0 100
rw 13 0 100

*Voltage source
vin 1 0 dc 5

*dc analysis 
.dc vin 0 10 0.01

.control
run

*plot the graphs required
plot i(v1) vs v(1,2) i(vr) vs v(1,3) i(vb) vs v(1,4) i(vy) vs v(1,5) i(vg) vs v(1,6) i(vw) vs v(1,7)

.endc
.end

