Lab3 Question1
.include Diode_1N914.txt
.include red_5mm.txt
.include green_5mm.txt
.include blue_5mm.txt
.include yellow_5mm.txt
.include white_5mm.txt

*defining the diode
d1 1 2 1N914
dr 1 3 RED
db 1 4 BLUE
dy 1 5 YELLOW
dg 1 6 GREEN
dw 1 7 WHITE

*Current sources for measuring current across diode
v1 2 0 dc 0 ac 0
vr 3 0 dc 0 ac 0
vb 4 0 dc 0 ac 0
vy 5 0 dc 0 ac 0
vg 6 0 dc 0 ac 0
vw 7 0 dc 0 ac 0

*Voltage source
vin 1 0 dc 5

*dc analysis 
.dc vin 0.001 10qui 0.01

.control
run

*plot the graphs required
plot ln(i(vr)) ln(i(vb)) ln(i(vg)) ln(i(vy)) ln(i(v1)) ln(i(vw))

.endc
.end

